`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:45:32 04/10/2018 
// Design Name: 
// Module Name:    frogger 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module frogger(ClkPort, vga_h_sync, vga_v_sync, vga_r, vga_g, vga_b, Sw0, Sw1, btnU, btnD, btnR, btnL,
	St_ce_bar, St_rp_bar, Mt_ce_bar, Mt_St_oe_bar, Mt_St_we_bar,
	An0, An1, An2, An3, Ca, Cb, Cc, Cd, Ce, Cf, Cg, Dp,
	LD0, LD1, LD2, LD3, LD4, LD5, LD6, LD7);
	input ClkPort, Sw0, btnU, btnD, btnR, btnL, Sw0, Sw1;
	output St_ce_bar, St_rp_bar, Mt_ce_bar, Mt_St_oe_bar, Mt_St_we_bar;
	output vga_h_sync, vga_v_sync, vga_r, vga_g, vga_b;
	output An0, An1, An2, An3, Ca, Cb, Cc, Cd, Ce, Cf, Cg, Dp;
	output LD0, LD1, LD2, LD3, LD4, LD5, LD6, LD7;
	reg vga_r, vga_g, vga_b;
	
	//////////////////////////////////////////////////////////////////////////////////////////
	
	/*  LOCAL SIGNALS */
	wire	reset, start, ClkPort, board_clk, clk, button_clk;
	
	BUF BUF1 (board_clk, ClkPort); 	
	BUF BUF2 (reset, Sw0);
	BUF BUF3 (start, Sw1);
	
	reg [27:0]	DIV_CLK;
	always @ (posedge board_clk, posedge reset)  
	begin : CLOCK_DIVIDER
      if (reset)
			DIV_CLK <= 0;
      else
			DIV_CLK <= DIV_CLK + 1'b1;
	end	

	assign	button_clk = DIV_CLK[18];
	assign	clk = DIV_CLK[1];
	assign 	{St_ce_bar, St_rp_bar, Mt_ce_bar, Mt_St_oe_bar, Mt_St_we_bar} = {5'b11111};
	
	wire inDisplayArea;
	wire [9:0] CounterX;
	wire [9:0] CounterY;

	hvsync_generator syncgen(.clk(clk), .reset(reset),.vga_h_sync(vga_h_sync), .vga_v_sync(vga_v_sync), .inDisplayArea(inDisplayArea), .CounterX(CounterX), .CounterY(CounterY));
	
	
	
	//counter counter1(.out(cnt1), .enable(1'b1), .clk(DIV_CLK[21]), .reset(1'b0));
	//counter counter2(.out(cnt2), .enable(1'b1), .clk(DIV_CLK[26]), .reset(1'b0));
	/////////////////////////////////////////////////////////////////
	///////////////		VGA control starts here		/////////////////
	/////////////////////////////////////////////////////////////////
	reg [9:0] position;
	reg [9:0] h_position;
	reg [9:0] cnt, cnt2, cnt3;
	
	always @(posedge DIV_CLK[21])
		begin
			if(reset)
				begin
					position<=500;
					h_position<=240;
				end
			else if(btnD && ~btnU)
				position<=position+2;
			else if(btnU && ~btnD)
				position<=position-2;
			else if(btnR && ~btnL)
				h_position<=h_position+2;
			else if(btnL && ~btnR)
				h_position<=h_position-2;
		end
	
	always @(posedge DIV_CLK[24])
		begin
			if(reset || (cnt>480))
				begin
					cnt<=0;
				end
			else
				cnt<=cnt+5;
		end
	always @(posedge DIV_CLK[23])
		begin
			if(reset || (cnt2>480))
				begin
					cnt2<=0;
				end
			else
				cnt2<=cnt2+5;
		end
	always @(posedge DIV_CLK[22])
		begin
			if(reset || (cnt3>480))
				begin
					cnt3<=0;
				end
			else
				cnt3<=cnt3+5;
		end
		
	wire frog = CounterY>=(position-10) && CounterY<=(position+10) && CounterX>=(h_position-10) && CounterX<=(h_position+10);
	//wire R = CounterX>(cnt) && CounterX<(50+cnt) && CounterY[5:3]==7;
	wire car1 = CounterX>(cnt) && CounterX<(50+cnt) && CounterY>30 && CounterY<50;
	wire car2 = CounterX>(cnt2) && CounterX<(50+cnt2) && CounterY>80 && CounterY<100;
	wire car3 = CounterX>(cnt3) && CounterX<(50+cnt3) && CounterY>140 && CounterY<160;
	wire car4 = CounterX>(cnt) && CounterX<(50+cnt) && CounterY>200 && CounterY<220;
	wire car5 = CounterX>(cnt2) && CounterX<(50+cnt2) && CounterY>300 && CounterY<320;
	
	wire hit_car1, hit_car2, hit_car3, hit_car4, hit_car5;
	assign hit_car1 = ( ((((position-10)>=30) && ((position-10)<=50)) || (((position+10)>=30) && ((position+10)<=50))) 
		&& ( (((h_position-10)>=(cnt)) && ((h_position-10)<=(50+cnt))) || (((h_position+10)>=(cnt)) && ((h_position+10)<=(50+cnt))) ) );
	
	assign hit = hit_car1;
	always @(posedge clk)
	begin
		vga_r <= (car1||car2||car3||car4||car5) & inDisplayArea & (state==ingame);
		vga_g <= frog & inDisplayArea & (state==ingame);
		vga_b <= vga_r & inDisplayArea & (state==ingame);
	end
	
	/////////////////////////////////////////////////////////////////
	//////////////  	  VGA control ends here 	 ///////////////////
	/////////////////////////////////////////////////////////////////
	
	reg[3:0] state;
	
	//reg[1:0] frogs = 2'b11;
	integer frogs = 3;
	// state declaration
   localparam  [1:0]
      newgame = 4'b0001,
      ingame    = 4'b0010,
      newlife = 4'b0100,
      done    = 4'b1000;
		
		assign ack = btnR&&(state==done);
		assign ack2 = btnL&&(state==done);
always @ (posedge clk, posedge reset)
	begin
		if(reset)
			begin
				if(ack2)
					state <= newgame;
				//frogs <= 3;
			end
		else
		begin
			case(state)
				newgame:
					begin
						state<=ingame;
						frogs<=3;
					end
				ingame:
					begin
						if(hit)
							frogs<=frogs-1;
							if(frogs==1)
								state<=done;
					end
				//newlife:
				
				done:
					begin
						if(ack)
							state<=newgame;
					end
			endcase			
		end
	end
	
	//OFL


/*		
	always @ (posedge Clk, posedge reset)
	begin
		if(reset)
			state <= QINIT;
		else
		begin
			case(state)
		
				QINIT:
					begin
					if({U,Z}==2'b10)
						state <= QG1GET;
					end
				QG1GET:
					if(~U)
						state <= QG1;
				QG1:
					if({U,Z}==2'b01)
						state <= QG10GET;
					else if(U)
						state <= QBAD;
				QG10GET:
					if(~Z)
						state <= QG10;
				QG10:
					if({U,Z}==2'b10)
						state <= QG101GET;
					else if(Z)
						state <= QBAD;
				QG101GET:
					if(~U)
						state <= QG101;
				QG101:
					if({U,Z}==2'b10)
						//state <= QG1011GET;
						state <= QG1011GET;
					else if(Z)
						state <= QBAD;
				QG1011GET:
					if(~U)
						state <= QG1011;
				QG1011:
					state <= QOPENING;
				QOPENING:
					if(TO)
						state <= QINIT;
				QBAD:
					if({U,Z}==2'b00)
						state <= QINIT;
			endcase			
		end
	end
	
	//OFL
	assign Unlock = QOPENING;
*/
		
	/////////////////////////////////////////////////////////////////
	//////////////  	  LD control starts here 	 ///////////////////
	/////////////////////////////////////////////////////////////////
	`define QI 			2'b00
	`define QGAME_1 	2'b01
	`define QGAME_2 	2'b10
	`define QDONE 		2'b11
	
	reg [3:0] p2_score;
	reg [3:0] p1_score;
	reg [1:0] sstate;
	wire LD0, LD1, LD2, LD3, LD4, LD5, LD6, LD7;
	
	assign LD0 = (p1_score == 4'b1010);
	assign LD1 = (p2_score == 4'b1010);
	
	assign LD2 = hit_car1;
	assign LD4 = reset;
	
	assign LD3 = (sstate == `QI);
	assign LD5 = (sstate == `QGAME_1);	
	assign LD6 = (sstate == `QGAME_2);
	assign LD7 = (sstate == `QDONE);
	
	/////////////////////////////////////////////////////////////////
	//////////////  	  LD control ends here 	 	////////////////////
	/////////////////////////////////////////////////////////////////
	
	/////////////////////////////////////////////////////////////////
	//////////////  	  SSD control starts here 	 ///////////////////
	/////////////////////////////////////////////////////////////////
	reg 	[3:0]	SSD;
	wire 	[3:0]	SSD0, SSD1, SSD2, SSD3;
	wire 	[1:0] ssdscan_clk;
	
	assign SSD3 = 4'b1111;
	assign SSD2 = 4'b1111;
	assign SSD1 = 4'b1111;
	assign SSD0 = position[3:0];
	
	// need a scan clk for the seven segment display 
	// 191Hz (50MHz / 2^18) works well
	assign ssdscan_clk = DIV_CLK[19:18];	
	assign An0	= !(~(ssdscan_clk[1]) && ~(ssdscan_clk[0]));  // when ssdscan_clk = 00
	assign An1	= !(~(ssdscan_clk[1]) &&  (ssdscan_clk[0]));  // when ssdscan_clk = 01
	assign An2	= !( (ssdscan_clk[1]) && ~(ssdscan_clk[0]));  // when ssdscan_clk = 10
	assign An3	= !( (ssdscan_clk[1]) &&  (ssdscan_clk[0]));  // when ssdscan_clk = 11
	
	always @ (ssdscan_clk, SSD0, SSD1, SSD2, SSD3)
	begin : SSD_SCAN_OUT
		case (ssdscan_clk) 
			2'b00:
					SSD = SSD0;
			2'b01:
					SSD = SSD1;
			2'b10:
					SSD = SSD2;
			2'b11:
					SSD = SSD3;
		endcase 
	end	

	// and finally convert SSD_num to ssd
	reg [6:0]  SSD_CATHODES;
	assign {Ca, Cb, Cc, Cd, Ce, Cf, Cg, Dp} = {SSD_CATHODES, 1'b1};
	// Following is Hex-to-SSD conversion
	always @ (SSD) 
	begin : HEX_TO_SSD
		case (SSD)		
			4'b1111: SSD_CATHODES = 7'b1111111 ; //Nothing 
			4'b0000: SSD_CATHODES = 7'b0000001 ; //0
			4'b0001: SSD_CATHODES = 7'b1001111 ; //1
			4'b0010: SSD_CATHODES = 7'b0010010 ; //2
			4'b0011: SSD_CATHODES = 7'b0000110 ; //3
			4'b0100: SSD_CATHODES = 7'b1001100 ; //4
			4'b0101: SSD_CATHODES = 7'b0100100 ; //5
			4'b0110: SSD_CATHODES = 7'b0100000 ; //6
			4'b0111: SSD_CATHODES = 7'b0001111 ; //7
			4'b1000: SSD_CATHODES = 7'b0000000 ; //8
			4'b1001: SSD_CATHODES = 7'b0000100 ; //9
			4'b1010: SSD_CATHODES = 7'b0001000 ; //10 or A
			default: SSD_CATHODES = 7'bXXXXXXX ; // default is not needed as we covered all cases
		endcase
	end
	
	/////////////////////////////////////////////////////////////////
	//////////////  	  SSD control ends here 	 ///////////////////
	/////////////////////////////////////////////////////////////////
endmodule